
//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Sun Apr  7 21:42:00 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_run_staller
// ------------------------------------------------------------------


module fir_run_staller (
  run_wen, input_rsci_wen_comp, output_rsci_wen_comp
);
  output run_wen;
  input input_rsci_wen_comp;
  input output_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = input_rsci_wen_comp & output_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_output_rsci_output_wait_dp
// ------------------------------------------------------------------


module fir_run_output_rsci_output_wait_dp (
  clk, rst, output_rsci_oswt, output_rsci_wen_comp, output_rsci_biwt, output_rsci_bdwt,
      output_rsci_bcwt
);
  input clk;
  input rst;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input output_rsci_biwt;
  input output_rsci_bdwt;
  output output_rsci_bcwt;
  reg output_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_wen_comp = (~ output_rsci_oswt) | output_rsci_biwt | output_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_bcwt <= 1'b0;
    end
    else begin
      output_rsci_bcwt <= ~((~(output_rsci_bcwt | output_rsci_biwt)) | output_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_output_rsci_output_wait_ctrl
// ------------------------------------------------------------------


module fir_run_output_rsci_output_wait_ctrl (
  run_wen, output_rsci_oswt, output_rsci_biwt, output_rsci_bdwt, output_rsci_bcwt,
      output_rsci_irdy, output_rsci_ivld_run_sct
);
  input run_wen;
  input output_rsci_oswt;
  output output_rsci_biwt;
  output output_rsci_bdwt;
  input output_rsci_bcwt;
  input output_rsci_irdy;
  output output_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire output_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_bdwt = output_rsci_oswt & run_wen;
  assign output_rsci_biwt = output_rsci_ogwt & output_rsci_irdy;
  assign output_rsci_ogwt = output_rsci_oswt & (~ output_rsci_bcwt);
  assign output_rsci_ivld_run_sct = output_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_input_rsci_input_wait_dp
// ------------------------------------------------------------------


module fir_run_input_rsci_input_wait_dp (
  clk, rst, input_rsci_oswt, input_rsci_wen_comp, input_rsci_idat_mxwt, input_rsci_biwt,
      input_rsci_bdwt, input_rsci_bcwt, input_rsci_idat
);
  input clk;
  input rst;
  input input_rsci_oswt;
  output input_rsci_wen_comp;
  output [7:0] input_rsci_idat_mxwt;
  input input_rsci_biwt;
  input input_rsci_bdwt;
  output input_rsci_bcwt;
  reg input_rsci_bcwt;
  input [7:0] input_rsci_idat;


  // Interconnect Declarations
  reg [7:0] input_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_rsci_wen_comp = (~ input_rsci_oswt) | input_rsci_biwt | input_rsci_bcwt;
  assign input_rsci_idat_mxwt = MUX_v_8_2_2(input_rsci_idat, input_rsci_idat_bfwt,
      input_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      input_rsci_bcwt <= 1'b0;
    end
    else begin
      input_rsci_bcwt <= ~((~(input_rsci_bcwt | input_rsci_biwt)) | input_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_rsci_idat_bfwt <= 8'b00000000;
    end
    else if ( input_rsci_biwt ) begin
      input_rsci_idat_bfwt <= input_rsci_idat;
    end
  end

  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_input_rsci_input_wait_ctrl
// ------------------------------------------------------------------


module fir_run_input_rsci_input_wait_ctrl (
  run_wen, input_rsci_oswt, input_rsci_biwt, input_rsci_bdwt, input_rsci_bcwt, input_rsci_irdy_run_sct,
      input_rsci_ivld
);
  input run_wen;
  input input_rsci_oswt;
  output input_rsci_biwt;
  output input_rsci_bdwt;
  input input_rsci_bcwt;
  output input_rsci_irdy_run_sct;
  input input_rsci_ivld;


  // Interconnect Declarations
  wire input_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_rsci_bdwt = input_rsci_oswt & run_wen;
  assign input_rsci_biwt = input_rsci_ogwt & input_rsci_ivld;
  assign input_rsci_ogwt = input_rsci_oswt & (~ input_rsci_bcwt);
  assign input_rsci_irdy_run_sct = input_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module decimator_run_run_fsm (
  clk, rst, run_wen, fsm_output
);
  input clk;
  input rst;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for decimator_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : decimator_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_staller
// ------------------------------------------------------------------


module decimator_run_staller (
  run_wen, din_rsci_wen_comp, dout_rsci_wen_comp
);
  output run_wen;
  input din_rsci_wen_comp;
  input dout_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = din_rsci_wen_comp & dout_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_dout_rsci_dout_wait_ctrl
// ------------------------------------------------------------------


module decimator_run_dout_rsci_dout_wait_ctrl (
  dout_rsci_iswt0, dout_rsci_biwt, dout_rsci_irdy
);
  input dout_rsci_iswt0;
  output dout_rsci_biwt;
  input dout_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_biwt = dout_rsci_iswt0 & dout_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_din_rsci_din_wait_ctrl
// ------------------------------------------------------------------


module decimator_run_din_rsci_din_wait_ctrl (
  din_rsci_iswt0, din_rsci_biwt, din_rsci_ivld
);
  input din_rsci_iswt0;
  output din_rsci_biwt;
  input din_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_biwt = din_rsci_iswt0 & din_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_output_rsci
// ------------------------------------------------------------------


module fir_run_output_rsci (
  clk, rst, output_rsc_dat, output_rsc_vld, output_rsc_rdy, run_wen, output_rsci_oswt,
      output_rsci_wen_comp, output_rsci_idat
);
  input clk;
  input rst;
  output [7:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input run_wen;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input [7:0] output_rsci_idat;


  // Interconnect Declarations
  wire output_rsci_biwt;
  wire output_rsci_bdwt;
  wire output_rsci_bcwt;
  wire output_rsci_irdy;
  wire output_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd8)) output_rsci (
      .irdy(output_rsci_irdy),
      .ivld(output_rsci_ivld_run_sct),
      .idat(output_rsci_idat),
      .rdy(output_rsc_rdy),
      .vld(output_rsc_vld),
      .dat(output_rsc_dat)
    );
  fir_run_output_rsci_output_wait_ctrl fir_run_output_rsci_output_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .output_rsci_oswt(output_rsci_oswt),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_bdwt(output_rsci_bdwt),
      .output_rsci_bcwt(output_rsci_bcwt),
      .output_rsci_irdy(output_rsci_irdy),
      .output_rsci_ivld_run_sct(output_rsci_ivld_run_sct)
    );
  fir_run_output_rsci_output_wait_dp fir_run_output_rsci_output_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .output_rsci_oswt(output_rsci_oswt),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_bdwt(output_rsci_bdwt),
      .output_rsci_bcwt(output_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_input_rsci
// ------------------------------------------------------------------


module fir_run_input_rsci (
  clk, rst, input_rsc_dat, input_rsc_vld, input_rsc_rdy, run_wen, input_rsci_oswt,
      input_rsci_wen_comp, input_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [7:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input run_wen;
  input input_rsci_oswt;
  output input_rsci_wen_comp;
  output [7:0] input_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_rsci_biwt;
  wire input_rsci_bdwt;
  wire input_rsci_bcwt;
  wire input_rsci_irdy_run_sct;
  wire input_rsci_ivld;
  wire [7:0] input_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd8)) input_rsci (
      .rdy(input_rsc_rdy),
      .vld(input_rsc_vld),
      .dat(input_rsc_dat),
      .irdy(input_rsci_irdy_run_sct),
      .ivld(input_rsci_ivld),
      .idat(input_rsci_idat)
    );
  fir_run_input_rsci_input_wait_ctrl fir_run_input_rsci_input_wait_ctrl_inst (
      .run_wen(run_wen),
      .input_rsci_oswt(input_rsci_oswt),
      .input_rsci_biwt(input_rsci_biwt),
      .input_rsci_bdwt(input_rsci_bdwt),
      .input_rsci_bcwt(input_rsci_bcwt),
      .input_rsci_irdy_run_sct(input_rsci_irdy_run_sct),
      .input_rsci_ivld(input_rsci_ivld)
    );
  fir_run_input_rsci_input_wait_dp fir_run_input_rsci_input_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .input_rsci_oswt(input_rsci_oswt),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .input_rsci_idat_mxwt(input_rsci_idat_mxwt),
      .input_rsci_biwt(input_rsci_biwt),
      .input_rsci_bdwt(input_rsci_bdwt),
      .input_rsci_bcwt(input_rsci_bcwt),
      .input_rsci_idat(input_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_dout_rsci
// ------------------------------------------------------------------


module decimator_run_dout_rsci (
  dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, dout_rsci_oswt, dout_rsci_wen_comp, dout_rsci_idat
);
  output [7:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input [7:0] dout_rsci_idat;


  // Interconnect Declarations
  wire dout_rsci_biwt;
  wire dout_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd6),
  .width(32'sd8)) dout_rsci (
      .irdy(dout_rsci_irdy),
      .ivld(dout_rsci_oswt),
      .idat(dout_rsci_idat),
      .rdy(dout_rsc_rdy),
      .vld(dout_rsc_vld),
      .dat(dout_rsc_dat)
    );
  decimator_run_dout_rsci_dout_wait_ctrl decimator_run_dout_rsci_dout_wait_ctrl_inst
      (
      .dout_rsci_iswt0(dout_rsci_oswt),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_irdy(dout_rsci_irdy)
    );
  assign dout_rsci_wen_comp = (~ dout_rsci_oswt) | dout_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_din_rsci
// ------------------------------------------------------------------


module decimator_run_din_rsci (
  din_rsc_dat, din_rsc_vld, din_rsc_rdy, din_rsci_oswt, din_rsci_wen_comp, din_rsci_idat_mxwt
);
  input [7:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [7:0] din_rsci_idat_mxwt;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_ivld;
  wire [7:0] din_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd5),
  .width(32'sd8)) din_rsci (
      .rdy(din_rsc_rdy),
      .vld(din_rsc_vld),
      .dat(din_rsc_dat),
      .irdy(din_rsci_oswt),
      .ivld(din_rsci_ivld),
      .idat(din_rsci_idat)
    );
  decimator_run_din_rsci_din_wait_ctrl decimator_run_din_rsci_din_wait_ctrl_inst
      (
      .din_rsci_iswt0(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_ivld(din_rsci_ivld)
    );
  assign din_rsci_idat_mxwt = din_rsci_idat;
  assign din_rsci_wen_comp = (~ din_rsci_oswt) | din_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run
// ------------------------------------------------------------------


module fir_run (
  clk, rst, input_rsc_dat, input_rsc_vld, input_rsc_rdy, coeffs, output_rsc_dat,
      output_rsc_vld, output_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [63:0] coeffs;
  output [7:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire input_rsci_wen_comp;
  wire [7:0] input_rsci_idat_mxwt;
  wire output_rsci_wen_comp;
  reg [7:0] output_rsci_idat;
  wire [3:0] main_1_MAC_acc_2_tmp;
  wire [4:0] nl_main_1_MAC_acc_2_tmp;
  wire [3:0] main_1_SHIFT_acc_1_tmp;
  wire [4:0] nl_main_1_SHIFT_acc_1_tmp;
  wire [3:0] main_2_MAC_acc_2_tmp;
  wire [4:0] nl_main_2_MAC_acc_2_tmp;
  wire [3:0] main_2_SHIFT_acc_1_tmp;
  wire [4:0] nl_main_2_SHIFT_acc_1_tmp;
  wire or_dcpl_7;
  wire nor_tmp_1;
  wire and_dcpl_5;
  wire and_dcpl_11;
  wire or_dcpl_14;
  wire or_dcpl_15;
  wire or_dcpl_16;
  wire or_dcpl_17;
  wire or_dcpl_18;
  wire or_dcpl_19;
  wire or_dcpl_20;
  wire or_dcpl_21;
  wire or_dcpl_22;
  wire or_dcpl_23;
  wire or_dcpl_24;
  wire or_dcpl_25;
  wire or_dcpl_26;
  wire and_dcpl_37;
  wire or_dcpl_32;
  reg lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1;
  reg lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0;
  reg [2:0] SHIFT_i_3_0_1_lpi_1_2_0;
  wire lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1_1;
  wire SHIFT_SHIFT_nor_4_ssc_1;
  wire SHIFT_and_17_cse_1;
  wire SHIFT_equal_tmp_2;
  wire [2:0] SHIFT_i_3_0_1_lpi_1_dfm_2_0_mx0w0;
  wire lfst_exit_main_2_SHIFT_lpi_1_dfm_1_1;
  wire lfst_exit_main_2_SHIFT_lpi_1_dfm_0_1;
  reg exitL_exit_main_2_SHIFT_sva;
  reg lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_0;
  reg lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_1;
  reg SHIFT_and_1_svs_st_1;
  reg main_stage_0_2;
  reg SHIFT_unequal_tmp_1_1;
  reg SHIFT_equal_tmp_1_1;
  reg SHIFT_and_1_svs;
  reg reg_output_rsci_oswt_cse;
  reg reg_input_rsci_oswt_cse;
  wire and_47_cse;
  wire and_48_cse;
  wire or_10_cse;
  wire mux_6_cse;
  wire MAC_nor_m1c;
  wire [7:0] z_out;
  reg [18:0] temp_1_lpi_1;
  reg [18:0] temp_lpi_1;
  reg [7:0] regs_3_sva;
  reg [7:0] regs_4_sva;
  reg [7:0] regs_2_sva;
  reg [7:0] regs_5_sva;
  reg [7:0] regs_1_sva;
  reg [7:0] regs_6_sva;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_7_sva;
  reg [7:0] regs_7_sva_dfm_1_1;
  reg [7:0] regs_6_sva_dfm_1_1;
  reg [7:0] regs_5_sva_dfm_1_1;
  reg [7:0] regs_4_sva_dfm_1_1;
  reg [7:0] regs_3_sva_dfm_1_1;
  reg [7:0] regs_2_sva_dfm_1_1;
  reg [7:0] regs_1_sva_dfm_1_1;
  reg SHIFT_asn_1_itm_1;
  reg [7:0] MAC_mux_itm_1;
  reg [2:0] main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1;
  reg [2:0] MAC_i_3_0_1_lpi_1_2_0;
  wire output_rsci_idat_mx0c1;
  wire [18:0] temp_1_sva_2;
  wire [19:0] nl_temp_1_sva_2;
  wire [18:0] temp_1_lpi_1_dfm_1;
  wire [2:0] MAC_i_3_0_1_lpi_1_dfm_2_0_mx0w0;
  wire [7:0] regs_0_sva_mx0;
  wire [18:0] temp_sva_2;
  wire [19:0] nl_temp_sva_2;
  wire SHIFT_and_1_svs_mx1c1;
  wire [7:0] MAC_mux_5;
  wire MAC_i_and_cse;
  wire MAC_and_9_cse;
  wire SHIFT_i_and_cse;
  wire or_49_cse;

  wire[18:0] SHIFT_SHIFT_and_4_nl;
  wire SHIFT_not_13_nl;
  wire SHIFT_SHIFT_or_nl;
  wire[2:0] SHIFT_SHIFT_SHIFT_or_nl;
  wire reg_regs_5_rgt_nl;
  wire SHIFT_regs_nor_nl;
  wire reg_regs_1_rgt_nl;
  wire SHIFT_regs_nor_1_nl;
  wire reg_regs_6_rgt_nl;
  wire SHIFT_regs_nor_2_nl;
  wire reg_regs_2_rgt_nl;
  wire SHIFT_regs_nor_3_nl;
  wire reg_regs_7_rgt_nl;
  wire mux_3_nl;
  wire mux_2_nl;
  wire or_13_nl;
  wire or_11_nl;
  wire reg_regs_3_rgt_nl;
  wire SHIFT_regs_nor_4_nl;
  wire reg_regs_4_rgt_nl;
  wire SHIFT_regs_nor_5_nl;
  wire[2:0] SHIFT_SHIFT_SHIFT_or_1_nl;
  wire[15:0] main_1_MAC_mul_nl;
  wire signed [15:0] nl_main_1_MAC_mul_sgnd;
  wire SHIFT_not_12_nl;
  wire SHIFT_and_nl;
  wire[15:0] main_2_MAC_mul_nl;
  wire[7:0] MAC_mux_2_nl;
  wire signed [15:0] nl_main_2_MAC_mul_sgnd;
  wire SHIFT_mux_26_nl;
  wire MAC_and_nl;
  wire MAC_and_1_nl;
  wire MAC_and_2_nl;
  wire MAC_and_3_nl;
  wire MAC_and_4_nl;
  wire MAC_and_5_nl;
  wire MAC_and_6_nl;
  wire MAC_and_7_nl;
  wire MAC_and_8_nl;
  wire[2:0] SHIFT_else_mux_15_nl;
  wire and_64_nl;

  // Interconnect Declarations for Component Instantiations 
  fir_run_input_rsci fir_run_input_rsci_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .run_wen(run_wen),
      .input_rsci_oswt(reg_input_rsci_oswt_cse),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .input_rsci_idat_mxwt(input_rsci_idat_mxwt)
    );
  fir_run_output_rsci fir_run_output_rsci_inst (
      .clk(clk),
      .rst(rst),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .run_wen(run_wen),
      .output_rsci_oswt(reg_output_rsci_oswt_cse),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_idat(output_rsci_idat)
    );
  fir_run_staller fir_run_staller_inst (
      .run_wen(run_wen),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .output_rsci_wen_comp(output_rsci_wen_comp)
    );
  assign MAC_and_9_cse = run_wen & or_10_cse;
  assign MAC_i_and_cse = run_wen & ((~ lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0) | exitL_exit_main_2_SHIFT_sva
      | (~ lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1));
  assign or_49_cse = (SHIFT_i_3_0_1_lpi_1_2_0!=3'b000);
  assign SHIFT_i_and_cse = run_wen & (or_dcpl_7 | lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0
      | or_10_cse);
  assign and_47_cse = (main_2_MAC_acc_2_tmp[3]) & (main_2_SHIFT_acc_1_tmp[3]);
  assign and_48_cse = (main_1_MAC_acc_2_tmp[3]) & (main_1_SHIFT_acc_1_tmp[3]);
  assign or_10_cse = (~ lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1) | exitL_exit_main_2_SHIFT_sva;
  assign mux_6_cse = MUX_s_1_2_2((~ lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0), and_48_cse,
      or_10_cse);
  assign nl_main_1_MAC_mul_sgnd = $signed(MAC_mux_itm_1) * $signed(MAC_mux_5);
  assign main_1_MAC_mul_nl = $unsigned(nl_main_1_MAC_mul_sgnd);
  assign nl_temp_1_sva_2 = temp_1_lpi_1_dfm_1 + conv_s2s_16_19(main_1_MAC_mul_nl);
  assign temp_1_sva_2 = nl_temp_1_sva_2[18:0];
  assign SHIFT_not_12_nl = ~ SHIFT_asn_1_itm_1;
  assign temp_1_lpi_1_dfm_1 = MUX_v_19_2_2(19'b0000000000000000000, temp_1_lpi_1,
      SHIFT_not_12_nl);
  assign MAC_i_3_0_1_lpi_1_dfm_2_0_mx0w0 = MUX_v_3_2_2(MAC_i_3_0_1_lpi_1_2_0, 3'b111,
      exitL_exit_main_2_SHIFT_sva);
  assign SHIFT_and_nl = (~ SHIFT_unequal_tmp_1_1) & main_stage_0_2;
  assign regs_0_sva_mx0 = MUX_v_8_2_2(regs_0_sva, input_rsci_idat_mxwt, SHIFT_and_nl);
  assign SHIFT_i_3_0_1_lpi_1_dfm_2_0_mx0w0 = MUX_v_3_2_2(SHIFT_i_3_0_1_lpi_1_2_0,
      3'b111, exitL_exit_main_2_SHIFT_sva);
  assign MAC_mux_2_nl = MUX_v_8_8_2((coeffs[7:0]), (coeffs[15:8]), (coeffs[23:16]),
      (coeffs[31:24]), (coeffs[39:32]), (coeffs[47:40]), (coeffs[55:48]), (coeffs[63:56]),
      main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1);
  assign nl_main_2_MAC_mul_sgnd = $signed(MAC_mux_2_nl) * $signed(MAC_mux_5);
  assign main_2_MAC_mul_nl = $unsigned(nl_main_2_MAC_mul_sgnd);
  assign nl_temp_sva_2 = temp_lpi_1 + conv_s2s_16_19(main_2_MAC_mul_nl);
  assign temp_sva_2 = nl_temp_sva_2[18:0];
  assign lfst_exit_main_2_SHIFT_lpi_1_dfm_1_1 = lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1
      & (~ exitL_exit_main_2_SHIFT_sva);
  assign lfst_exit_main_2_SHIFT_lpi_1_dfm_0_1 = lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0
      & (~ exitL_exit_main_2_SHIFT_sva);
  assign SHIFT_mux_26_nl = MUX_s_1_2_2(and_47_cse, SHIFT_and_1_svs, or_dcpl_32);
  assign lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1_1 = (~(SHIFT_mux_26_nl | SHIFT_SHIFT_nor_4_ssc_1))
      | SHIFT_and_17_cse_1;
  assign SHIFT_SHIFT_nor_4_ssc_1 = ~(and_48_cse | SHIFT_equal_tmp_2);
  assign SHIFT_equal_tmp_2 = lfst_exit_main_2_SHIFT_lpi_1_dfm_1_1 & (~ lfst_exit_main_2_SHIFT_lpi_1_dfm_0_1);
  assign nl_main_1_SHIFT_acc_1_tmp = conv_u2s_3_4(SHIFT_i_3_0_1_lpi_1_dfm_2_0_mx0w0)
      + 4'b1111;
  assign main_1_SHIFT_acc_1_tmp = nl_main_1_SHIFT_acc_1_tmp[3:0];
  assign SHIFT_and_17_cse_1 = and_48_cse & (~ SHIFT_equal_tmp_2);
  assign nl_main_1_MAC_acc_2_tmp = conv_u2s_3_4(MAC_i_3_0_1_lpi_1_dfm_2_0_mx0w0)
      + 4'b1111;
  assign main_1_MAC_acc_2_tmp = nl_main_1_MAC_acc_2_tmp[3:0];
  assign nl_main_2_SHIFT_acc_1_tmp = conv_u2s_3_4(SHIFT_i_3_0_1_lpi_1_2_0) + 4'b1111;
  assign main_2_SHIFT_acc_1_tmp = nl_main_2_SHIFT_acc_1_tmp[3:0];
  assign nl_main_2_MAC_acc_2_tmp = conv_u2s_3_4(MAC_i_3_0_1_lpi_1_2_0) + 4'b1111;
  assign main_2_MAC_acc_2_tmp = nl_main_2_MAC_acc_2_tmp[3:0];
  assign MAC_nor_m1c = ~((main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1!=3'b000));
  assign MAC_and_nl = (~ SHIFT_unequal_tmp_1_1) & MAC_nor_m1c;
  assign MAC_and_1_nl = SHIFT_unequal_tmp_1_1 & MAC_nor_m1c;
  assign MAC_and_2_nl = (main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1==3'b001);
  assign MAC_and_3_nl = (main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1==3'b010);
  assign MAC_and_4_nl = (main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1==3'b011);
  assign MAC_and_5_nl = (main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1==3'b100);
  assign MAC_and_6_nl = (main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1==3'b101);
  assign MAC_and_7_nl = (main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1==3'b110);
  assign MAC_and_8_nl = (main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1==3'b111);
  assign MAC_mux_5 = MUX1HOT_v_8_9_2(input_rsci_idat_mxwt, regs_0_sva, regs_1_sva_dfm_1_1,
      regs_2_sva_dfm_1_1, regs_3_sva_dfm_1_1, regs_4_sva_dfm_1_1, regs_5_sva_dfm_1_1,
      regs_6_sva_dfm_1_1, regs_7_sva_dfm_1_1, {MAC_and_nl , MAC_and_1_nl , MAC_and_2_nl
      , MAC_and_3_nl , MAC_and_4_nl , MAC_and_5_nl , MAC_and_6_nl , MAC_and_7_nl
      , MAC_and_8_nl});
  assign or_dcpl_7 = ~((main_2_SHIFT_acc_1_tmp[3]) & (main_2_MAC_acc_2_tmp[3]));
  assign nor_tmp_1 = (main_1_SHIFT_acc_1_tmp[2:0]==3'b111);
  assign and_dcpl_5 = main_stage_0_2 & SHIFT_and_1_svs_st_1;
  assign and_dcpl_11 = main_stage_0_2 & (~ SHIFT_equal_tmp_1_1);
  assign or_dcpl_14 = (SHIFT_i_3_0_1_lpi_1_2_0[2]) | exitL_exit_main_2_SHIFT_sva;
  assign or_dcpl_15 = (SHIFT_i_3_0_1_lpi_1_2_0[1:0]!=2'b01);
  assign or_dcpl_16 = or_dcpl_15 | or_dcpl_14;
  assign or_dcpl_17 = (SHIFT_i_3_0_1_lpi_1_2_0[1:0]!=2'b10);
  assign or_dcpl_18 = or_dcpl_17 | or_dcpl_14;
  assign or_dcpl_19 = ~((SHIFT_i_3_0_1_lpi_1_2_0[1:0]==2'b11));
  assign or_dcpl_20 = or_dcpl_19 | or_dcpl_14;
  assign or_dcpl_21 = (~ (SHIFT_i_3_0_1_lpi_1_2_0[2])) | exitL_exit_main_2_SHIFT_sva;
  assign or_dcpl_22 = (SHIFT_i_3_0_1_lpi_1_2_0[1:0]!=2'b00);
  assign or_dcpl_23 = or_dcpl_22 | or_dcpl_21;
  assign or_dcpl_24 = or_dcpl_15 | or_dcpl_21;
  assign or_dcpl_25 = or_dcpl_17 | or_dcpl_21;
  assign or_dcpl_26 = or_dcpl_19 | (~ (SHIFT_i_3_0_1_lpi_1_2_0[2]));
  assign and_dcpl_37 = or_dcpl_26 & (~ exitL_exit_main_2_SHIFT_sva);
  assign or_dcpl_32 = lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0 | exitL_exit_main_2_SHIFT_sva
      | (~ lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1);
  assign output_rsci_idat_mx0c1 = and_dcpl_5 & (~ lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_0)
      & lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_1;
  assign SHIFT_and_1_svs_mx1c1 = and_48_cse & or_10_cse;
  always @(posedge clk) begin
    if ( rst ) begin
      reg_output_rsci_oswt_cse <= 1'b0;
      lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_1 <= 1'b0;
      lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_0 <= 1'b0;
      reg_input_rsci_oswt_cse <= 1'b0;
      lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1 <= 1'b0;
      exitL_exit_main_2_SHIFT_sva <= 1'b1;
      lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      SHIFT_equal_tmp_1_1 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_output_rsci_oswt_cse <= ~((~(main_stage_0_2 & SHIFT_and_1_svs_st_1)) |
          (lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_0 & lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_1));
      lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_1 <= lfst_exit_main_2_SHIFT_lpi_1_dfm_1_1;
      lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_0 <= lfst_exit_main_2_SHIFT_lpi_1_dfm_0_1;
      reg_input_rsci_oswt_cse <= ~(or_dcpl_22 | (SHIFT_i_3_0_1_lpi_1_2_0[2]) | (lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0
          & lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1) | exitL_exit_main_2_SHIFT_sva);
      lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1 <= lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1_1;
      exitL_exit_main_2_SHIFT_sva <= ~(lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1_1 | SHIFT_SHIFT_nor_4_ssc_1);
      lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0 <= SHIFT_SHIFT_nor_4_ssc_1;
      main_stage_0_2 <= 1'b1;
      SHIFT_equal_tmp_1_1 <= SHIFT_equal_tmp_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat <= 8'b00000000;
    end
    else if ( run_wen & ((and_dcpl_5 & (~ lfst_exit_main_2_SHIFT_lpi_1_dfm_st_1_1))
        | output_rsci_idat_mx0c1) ) begin
      output_rsci_idat <= MUX_v_8_2_2((temp_1_sva_2[18:11]), (temp_sva_2[18:11]),
          output_rsci_idat_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_mux_itm_1 <= 8'b00000000;
      SHIFT_asn_1_itm_1 <= 1'b0;
    end
    else if ( MAC_and_9_cse ) begin
      MAC_mux_itm_1 <= MUX_v_8_8_2((coeffs[7:0]), (coeffs[15:8]), (coeffs[23:16]),
          (coeffs[31:24]), (coeffs[39:32]), (coeffs[47:40]), (coeffs[55:48]), (coeffs[63:56]),
          MAC_i_3_0_1_lpi_1_dfm_2_0_mx0w0);
      SHIFT_asn_1_itm_1 <= exitL_exit_main_2_SHIFT_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1 <= 3'b000;
      SHIFT_and_1_svs_st_1 <= 1'b0;
      regs_1_sva_dfm_1_1 <= 8'b00000000;
      regs_2_sva_dfm_1_1 <= 8'b00000000;
      regs_3_sva_dfm_1_1 <= 8'b00000000;
      regs_4_sva_dfm_1_1 <= 8'b00000000;
      regs_5_sva_dfm_1_1 <= 8'b00000000;
      regs_6_sva_dfm_1_1 <= 8'b00000000;
      regs_7_sva_dfm_1_1 <= 8'b00000000;
      SHIFT_unequal_tmp_1_1 <= 1'b0;
    end
    else if ( MAC_i_and_cse ) begin
      main_1_MAC_i_slc_MAC_i_3_0_2_0_itm_1 <= MUX_v_3_2_2(MAC_i_3_0_1_lpi_1_dfm_2_0_mx0w0,
          MAC_i_3_0_1_lpi_1_2_0, lfst_exit_main_2_SHIFT_lpi_1_dfm_1_1);
      SHIFT_and_1_svs_st_1 <= MUX_s_1_2_2(and_47_cse, and_48_cse, or_10_cse);
      regs_1_sva_dfm_1_1 <= MUX_v_8_2_2(z_out, regs_1_sva, or_dcpl_16);
      regs_2_sva_dfm_1_1 <= MUX_v_8_2_2(z_out, regs_2_sva, or_dcpl_18);
      regs_3_sva_dfm_1_1 <= MUX_v_8_2_2(z_out, regs_3_sva, or_dcpl_20);
      regs_4_sva_dfm_1_1 <= MUX_v_8_2_2(z_out, regs_4_sva, or_dcpl_23);
      regs_5_sva_dfm_1_1 <= MUX_v_8_2_2(z_out, regs_5_sva, or_dcpl_24);
      regs_6_sva_dfm_1_1 <= MUX_v_8_2_2(z_out, regs_6_sva, or_dcpl_25);
      regs_7_sva_dfm_1_1 <= MUX_v_8_2_2(z_out, regs_7_sva, and_dcpl_37);
      SHIFT_unequal_tmp_1_1 <= MUX_s_1_2_2(or_49_cse, SHIFT_SHIFT_or_nl, or_10_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_0_sva <= 8'b00000000;
    end
    else if ( ((or_49_cse & (~(lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1 & lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0)))
        | exitL_exit_main_2_SHIFT_sva) & run_wen & (~ SHIFT_unequal_tmp_1_1) & main_stage_0_2
        ) begin
      regs_0_sva <= regs_0_sva_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      temp_lpi_1 <= 19'b0000000000000000000;
    end
    else if ( lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1 & (~ exitL_exit_main_2_SHIFT_sva)
        & (SHIFT_and_1_svs | SHIFT_equal_tmp_1_1) & (~ lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0)
        & main_stage_0_2 & run_wen ) begin
      temp_lpi_1 <= MUX_v_19_2_2(temp_sva_2, SHIFT_SHIFT_and_4_nl, and_dcpl_11);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      temp_1_lpi_1 <= 19'b0000000000000000000;
    end
    else if ( run_wen & main_stage_0_2 & (~ lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1)
        & (~((~(SHIFT_asn_1_itm_1 | (~ SHIFT_equal_tmp_1_1))) | exitL_exit_main_2_SHIFT_sva))
        ) begin
      temp_1_lpi_1 <= MUX_v_19_2_2(temp_1_lpi_1_dfm_1, temp_1_sva_2, and_dcpl_11);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      SHIFT_i_3_0_1_lpi_1_2_0 <= 3'b000;
      MAC_i_3_0_1_lpi_1_2_0 <= 3'b000;
    end
    else if ( SHIFT_i_and_cse ) begin
      SHIFT_i_3_0_1_lpi_1_2_0 <= MUX_v_3_2_2((main_1_SHIFT_acc_1_tmp[2:0]), SHIFT_SHIFT_SHIFT_or_nl,
          mux_6_cse);
      MAC_i_3_0_1_lpi_1_2_0 <= MUX_v_3_2_2((main_1_MAC_acc_2_tmp[2:0]), SHIFT_SHIFT_SHIFT_or_1_nl,
          mux_6_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_5_sva <= 8'b00000000;
    end
    else if ( run_wen & reg_regs_5_rgt_nl ) begin
      regs_5_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_1_sva <= 8'b00000000;
    end
    else if ( run_wen & reg_regs_1_rgt_nl ) begin
      regs_1_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_6_sva <= 8'b00000000;
    end
    else if ( run_wen & reg_regs_6_rgt_nl ) begin
      regs_6_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_2_sva <= 8'b00000000;
    end
    else if ( run_wen & reg_regs_2_rgt_nl ) begin
      regs_2_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_7_sva <= 8'b00000000;
    end
    else if ( ~((~ run_wen) | reg_regs_7_rgt_nl | mux_3_nl) ) begin
      regs_7_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_3_sva <= 8'b00000000;
    end
    else if ( run_wen & reg_regs_3_rgt_nl ) begin
      regs_3_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_4_sva <= 8'b00000000;
    end
    else if ( run_wen & reg_regs_4_rgt_nl ) begin
      regs_4_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      SHIFT_and_1_svs <= 1'b0;
    end
    else if ( run_wen & (((~(lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0 | exitL_exit_main_2_SHIFT_sva))
        & lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1) | SHIFT_and_1_svs_mx1c1) & ((~ or_dcpl_7)
        | or_10_cse) ) begin
      SHIFT_and_1_svs <= MUX_s_1_2_2(and_47_cse, and_48_cse, SHIFT_and_1_svs_mx1c1);
    end
  end
  assign SHIFT_SHIFT_or_nl = (SHIFT_i_3_0_1_lpi_1_dfm_2_0_mx0w0!=3'b000);
  assign SHIFT_not_13_nl = ~ SHIFT_and_1_svs;
  assign SHIFT_SHIFT_and_4_nl = MUX_v_19_2_2(19'b0000000000000000000, temp_lpi_1,
      SHIFT_not_13_nl);
  assign SHIFT_SHIFT_SHIFT_or_nl = MUX_v_3_2_2((main_2_SHIFT_acc_1_tmp[2:0]), 3'b111,
      SHIFT_and_17_cse_1);
  assign SHIFT_SHIFT_SHIFT_or_1_nl = MUX_v_3_2_2((main_2_MAC_acc_2_tmp[2:0]), 3'b111,
      SHIFT_and_17_cse_1);
  assign SHIFT_regs_nor_nl = ~(or_dcpl_15 | (~ (SHIFT_i_3_0_1_lpi_1_2_0[2])));
  assign reg_regs_5_rgt_nl = MUX_s_1_2_2(SHIFT_regs_nor_nl, (~ or_dcpl_24), or_dcpl_32);
  assign SHIFT_regs_nor_1_nl = ~(or_dcpl_15 | (SHIFT_i_3_0_1_lpi_1_2_0[2]));
  assign reg_regs_1_rgt_nl = MUX_s_1_2_2(SHIFT_regs_nor_1_nl, (~ or_dcpl_16), or_dcpl_32);
  assign SHIFT_regs_nor_2_nl = ~(or_dcpl_17 | (~ (SHIFT_i_3_0_1_lpi_1_2_0[2])));
  assign reg_regs_6_rgt_nl = MUX_s_1_2_2(SHIFT_regs_nor_2_nl, (~ or_dcpl_25), or_dcpl_32);
  assign SHIFT_regs_nor_3_nl = ~(or_dcpl_17 | (SHIFT_i_3_0_1_lpi_1_2_0[2]));
  assign reg_regs_2_rgt_nl = MUX_s_1_2_2(SHIFT_regs_nor_3_nl, (~ or_dcpl_18), or_dcpl_32);
  assign reg_regs_7_rgt_nl = MUX_s_1_2_2(or_dcpl_26, and_dcpl_37, or_dcpl_32);
  assign or_13_nl = ((main_2_SHIFT_acc_1_tmp[2:0]==3'b111)) | and_47_cse;
  assign mux_2_nl = MUX_s_1_2_2(or_13_nl, nor_tmp_1, lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0);
  assign or_11_nl = and_48_cse | nor_tmp_1;
  assign mux_3_nl = MUX_s_1_2_2(mux_2_nl, or_11_nl, or_10_cse);
  assign SHIFT_regs_nor_4_nl = ~(or_dcpl_19 | (SHIFT_i_3_0_1_lpi_1_2_0[2]));
  assign reg_regs_3_rgt_nl = MUX_s_1_2_2(SHIFT_regs_nor_4_nl, (~ or_dcpl_20), or_dcpl_32);
  assign SHIFT_regs_nor_5_nl = ~(or_dcpl_22 | (~ (SHIFT_i_3_0_1_lpi_1_2_0[2])));
  assign reg_regs_4_rgt_nl = MUX_s_1_2_2(SHIFT_regs_nor_5_nl, (~ or_dcpl_23), or_dcpl_32);
  assign and_64_nl = lfst_exit_main_2_SHIFT_lpi_1_dfm_3_1 & (~ exitL_exit_main_2_SHIFT_sva)
      & (~ lfst_exit_main_2_SHIFT_lpi_1_dfm_3_0);
  assign SHIFT_else_mux_15_nl = MUX_v_3_2_2(SHIFT_i_3_0_1_lpi_1_dfm_2_0_mx0w0, SHIFT_i_3_0_1_lpi_1_2_0,
      and_64_nl);
  assign z_out = MUX_v_8_8_2x0(regs_0_sva_mx0, regs_1_sva, regs_2_sva, regs_3_sva,
      regs_4_sva, regs_5_sva, regs_6_sva, SHIFT_else_mux_15_nl);

  function automatic [7:0] MUX1HOT_v_8_9_2;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [8:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    result = result | (input_8 & {8{sel[8]}});
    MUX1HOT_v_8_9_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [18:0] MUX_v_19_2_2;
    input [18:0] input_0;
    input [18:0] input_1;
    input  sel;
    reg [18:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_19_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2x0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2x0 = result;
  end
  endfunction


  function automatic [18:0] conv_s2s_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run
// ------------------------------------------------------------------


module decimator_run (
  clk, rst, din_rsc_dat, din_rsc_vld, din_rsc_rdy, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  output [7:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire din_rsci_wen_comp;
  wire [7:0] din_rsci_idat_mxwt;
  wire dout_rsci_wen_comp;
  reg [7:0] dout_rsci_idat;
  wire [2:0] fsm_output;
  wire equal_tmp;
  reg reg_dout_rsci_iswt0_cse;
  reg reg_din_rsci_iswt0_cse;
  reg [1:0] count_2_0_sva_1_0;
  wire [2:0] nl_count_2_0_sva_1_0;


  // Interconnect Declarations for Component Instantiations 
  decimator_run_din_rsci decimator_run_din_rsci_inst (
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .din_rsci_oswt(reg_din_rsci_iswt0_cse),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt)
    );
  decimator_run_dout_rsci decimator_run_dout_rsci_inst (
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .dout_rsci_oswt(reg_dout_rsci_iswt0_cse),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_idat(dout_rsci_idat)
    );
  decimator_run_staller decimator_run_staller_inst (
      .run_wen(run_wen),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .dout_rsci_wen_comp(dout_rsci_wen_comp)
    );
  decimator_run_run_fsm decimator_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign equal_tmp = ~((count_2_0_sva_1_0!=2'b00));
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_idat <= 8'b00000000;
    end
    else if ( run_wen & equal_tmp & (fsm_output[1]) ) begin
      dout_rsci_idat <= din_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_dout_rsci_iswt0_cse <= 1'b0;
      reg_din_rsci_iswt0_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_dout_rsci_iswt0_cse <= equal_tmp & (fsm_output[1]);
      reg_din_rsci_iswt0_cse <= ~ (fsm_output[1]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      count_2_0_sva_1_0 <= 2'b00;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      count_2_0_sva_1_0 <= nl_count_2_0_sva_1_0[1:0];
    end
  end
  assign nl_count_2_0_sva_1_0  = count_2_0_sva_1_0 + 2'b01;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, input_rsc_dat, input_rsc_vld, input_rsc_rdy, coeffs, output_rsc_dat,
      output_rsc_vld, output_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [63:0] coeffs;
  output [7:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  fir_run fir_run_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .coeffs(coeffs),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator
// ------------------------------------------------------------------


module decimator (
  clk, rst, din_rsc_dat, din_rsc_vld, din_rsc_rdy, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  output [7:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  decimator_run decimator_run_inst (
      .clk(clk),
      .rst(rst),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    top
// ------------------------------------------------------------------


module top (
  clk, rst, din_rsc_dat, din_rsc_vld, din_rsc_rdy, coeffs, dout_rsc_dat, dout_rsc_vld,
      dout_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input [63:0] coeffs;
  output [7:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;


  // Interconnect Declarations
  wire [7:0] output_rsc_dat_n_block0;
  wire [7:0] output_rsc_dat_n_block1;
  wire [7:0] dout_rsc_dat_n_block2;
  wire input_rsc_rdy_n_block0_bud;
  wire output_rsc_vld_n_block0_bud;
  wire input_rsc_rdy_n_block1_bud;
  wire output_rsc_vld_n_block1_bud;
  wire din_rsc_rdy_n_block2_bud;
  wire dout_rsc_vld_n_block2_bud;


  // Interconnect Declarations for Component Instantiations 
  fir block0 (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(din_rsc_dat),
      .input_rsc_vld(din_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy_n_block0_bud),
      .coeffs(coeffs),
      .output_rsc_dat(output_rsc_dat_n_block0),
      .output_rsc_vld(output_rsc_vld_n_block0_bud),
      .output_rsc_rdy(input_rsc_rdy_n_block1_bud)
    );
  fir block1 (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(output_rsc_dat_n_block0),
      .input_rsc_vld(output_rsc_vld_n_block0_bud),
      .input_rsc_rdy(input_rsc_rdy_n_block1_bud),
      .coeffs(coeffs),
      .output_rsc_dat(output_rsc_dat_n_block1),
      .output_rsc_vld(output_rsc_vld_n_block1_bud),
      .output_rsc_rdy(din_rsc_rdy_n_block2_bud)
    );
  decimator block2 (
      .clk(clk),
      .rst(rst),
      .din_rsc_dat(output_rsc_dat_n_block1),
      .din_rsc_vld(output_rsc_vld_n_block1_bud),
      .din_rsc_rdy(din_rsc_rdy_n_block2_bud),
      .dout_rsc_dat(dout_rsc_dat_n_block2),
      .dout_rsc_vld(dout_rsc_vld_n_block2_bud),
      .dout_rsc_rdy(dout_rsc_rdy)
    );
  assign din_rsc_rdy = input_rsc_rdy_n_block0_bud;
  assign dout_rsc_vld = dout_rsc_vld_n_block2_bud;
  assign dout_rsc_dat = dout_rsc_dat_n_block2;
endmodule



