
//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m111061545@ws41
//  Generated date: Sun Apr  7 21:44:27 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_run_run_fsm (
  clk, rst, run_wen, fsm_output
);
  input clk;
  input rst;
  input run_wen;
  output [9:0] fsm_output;
  reg [9:0] fsm_output;


  // FSM State Type Declaration for fir_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    main_C_3 = 4'd4,
    main_C_4 = 4'd5,
    main_C_5 = 4'd6,
    main_C_6 = 4'd7,
    main_C_7 = 4'd8,
    main_C_8 = 4'd9;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 10'b0000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 10'b0000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 10'b0000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 10'b0000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 10'b0000100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 10'b0001000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 10'b0010000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 10'b0100000000;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 10'b1000000000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 10'b0000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_staller
// ------------------------------------------------------------------


module fir_run_staller (
  run_wen, input_rsci_wen_comp, output_rsci_wen_comp
);
  output run_wen;
  input input_rsci_wen_comp;
  input output_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = input_rsci_wen_comp & output_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_output_rsci_output_wait_ctrl
// ------------------------------------------------------------------


module fir_run_output_rsci_output_wait_ctrl (
  output_rsci_iswt0, output_rsci_biwt, output_rsci_irdy
);
  input output_rsci_iswt0;
  output output_rsci_biwt;
  input output_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_biwt = output_rsci_iswt0 & output_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_input_rsci_input_wait_ctrl
// ------------------------------------------------------------------


module fir_run_input_rsci_input_wait_ctrl (
  input_rsci_iswt0, input_rsci_biwt, input_rsci_ivld
);
  input input_rsci_iswt0;
  output input_rsci_biwt;
  input input_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign input_rsci_biwt = input_rsci_iswt0 & input_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module decimator_run_run_fsm (
  clk, rst, run_wen, fsm_output
);
  input clk;
  input rst;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for decimator_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : decimator_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_staller
// ------------------------------------------------------------------


module decimator_run_staller (
  run_wen, din_rsci_wen_comp, dout_rsci_wen_comp
);
  output run_wen;
  input din_rsci_wen_comp;
  input dout_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = din_rsci_wen_comp & dout_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_dout_rsci_dout_wait_dp
// ------------------------------------------------------------------


module decimator_run_dout_rsci_dout_wait_dp (
  clk, rst, dout_rsci_oswt, dout_rsci_wen_comp, dout_rsci_biwt, dout_rsci_bdwt, dout_rsci_bcwt
);
  input clk;
  input rst;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input dout_rsci_biwt;
  input dout_rsci_bdwt;
  output dout_rsci_bcwt;
  reg dout_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_wen_comp = (~ dout_rsci_oswt) | dout_rsci_biwt | dout_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_bcwt <= 1'b0;
    end
    else begin
      dout_rsci_bcwt <= ~((~(dout_rsci_bcwt | dout_rsci_biwt)) | dout_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_dout_rsci_dout_wait_ctrl
// ------------------------------------------------------------------


module decimator_run_dout_rsci_dout_wait_ctrl (
  run_wen, dout_rsci_oswt, dout_rsci_biwt, dout_rsci_bdwt, dout_rsci_bcwt, dout_rsci_irdy,
      dout_rsci_ivld_run_sct
);
  input run_wen;
  input dout_rsci_oswt;
  output dout_rsci_biwt;
  output dout_rsci_bdwt;
  input dout_rsci_bcwt;
  input dout_rsci_irdy;
  output dout_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire dout_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_bdwt = dout_rsci_oswt & run_wen;
  assign dout_rsci_biwt = dout_rsci_ogwt & dout_rsci_irdy;
  assign dout_rsci_ogwt = dout_rsci_oswt & (~ dout_rsci_bcwt);
  assign dout_rsci_ivld_run_sct = dout_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_din_rsci_din_wait_dp
// ------------------------------------------------------------------


module decimator_run_din_rsci_din_wait_dp (
  clk, rst, din_rsci_oswt, din_rsci_wen_comp, din_rsci_idat_mxwt, din_rsci_biwt,
      din_rsci_bdwt, din_rsci_bcwt, din_rsci_idat
);
  input clk;
  input rst;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [7:0] din_rsci_idat_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  output din_rsci_bcwt;
  reg din_rsci_bcwt;
  input [7:0] din_rsci_idat;


  // Interconnect Declarations
  reg [7:0] din_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_wen_comp = (~ din_rsci_oswt) | din_rsci_biwt | din_rsci_bcwt;
  assign din_rsci_idat_mxwt = MUX_v_8_2_2(din_rsci_idat, din_rsci_idat_bfwt, din_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsci_bcwt <= 1'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsci_idat_bfwt <= 8'b00000000;
    end
    else if ( din_rsci_biwt ) begin
      din_rsci_idat_bfwt <= din_rsci_idat;
    end
  end

  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_din_rsci_din_wait_ctrl
// ------------------------------------------------------------------


module decimator_run_din_rsci_din_wait_ctrl (
  run_wen, din_rsci_oswt, din_rsci_biwt, din_rsci_bdwt, din_rsci_bcwt, din_rsci_irdy_run_sct,
      din_rsci_ivld
);
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  input din_rsci_bcwt;
  output din_rsci_irdy_run_sct;
  input din_rsci_ivld;


  // Interconnect Declarations
  wire din_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & run_wen;
  assign din_rsci_biwt = din_rsci_ogwt & din_rsci_ivld;
  assign din_rsci_ogwt = din_rsci_oswt & (~ din_rsci_bcwt);
  assign din_rsci_irdy_run_sct = din_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_output_rsci
// ------------------------------------------------------------------


module fir_run_output_rsci (
  output_rsc_dat, output_rsc_vld, output_rsc_rdy, output_rsci_oswt, output_rsci_wen_comp,
      output_rsci_idat
);
  output [7:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input [7:0] output_rsci_idat;


  // Interconnect Declarations
  wire output_rsci_biwt;
  wire output_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd8)) output_rsci (
      .irdy(output_rsci_irdy),
      .ivld(output_rsci_oswt),
      .idat(output_rsci_idat),
      .rdy(output_rsc_rdy),
      .vld(output_rsc_vld),
      .dat(output_rsc_dat)
    );
  fir_run_output_rsci_output_wait_ctrl fir_run_output_rsci_output_wait_ctrl_inst
      (
      .output_rsci_iswt0(output_rsci_oswt),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_irdy(output_rsci_irdy)
    );
  assign output_rsci_wen_comp = (~ output_rsci_oswt) | output_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run_input_rsci
// ------------------------------------------------------------------


module fir_run_input_rsci (
  input_rsc_dat, input_rsc_vld, input_rsc_rdy, input_rsci_oswt, input_rsci_wen_comp,
      input_rsci_idat_mxwt
);
  input [7:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input input_rsci_oswt;
  output input_rsci_wen_comp;
  output [7:0] input_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_rsci_biwt;
  wire input_rsci_ivld;
  wire [7:0] input_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd8)) input_rsci (
      .rdy(input_rsc_rdy),
      .vld(input_rsc_vld),
      .dat(input_rsc_dat),
      .irdy(input_rsci_oswt),
      .ivld(input_rsci_ivld),
      .idat(input_rsci_idat)
    );
  fir_run_input_rsci_input_wait_ctrl fir_run_input_rsci_input_wait_ctrl_inst (
      .input_rsci_iswt0(input_rsci_oswt),
      .input_rsci_biwt(input_rsci_biwt),
      .input_rsci_ivld(input_rsci_ivld)
    );
  assign input_rsci_idat_mxwt = input_rsci_idat;
  assign input_rsci_wen_comp = (~ input_rsci_oswt) | input_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_dout_rsci
// ------------------------------------------------------------------


module decimator_run_dout_rsci (
  clk, rst, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, run_wen, dout_rsci_oswt, dout_rsci_wen_comp,
      dout_rsci_idat
);
  input clk;
  input rst;
  output [7:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  input run_wen;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input [7:0] dout_rsci_idat;


  // Interconnect Declarations
  wire dout_rsci_biwt;
  wire dout_rsci_bdwt;
  wire dout_rsci_bcwt;
  wire dout_rsci_irdy;
  wire dout_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd6),
  .width(32'sd8)) dout_rsci (
      .irdy(dout_rsci_irdy),
      .ivld(dout_rsci_ivld_run_sct),
      .idat(dout_rsci_idat),
      .rdy(dout_rsc_rdy),
      .vld(dout_rsc_vld),
      .dat(dout_rsc_dat)
    );
  decimator_run_dout_rsci_dout_wait_ctrl decimator_run_dout_rsci_dout_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt),
      .dout_rsci_irdy(dout_rsci_irdy),
      .dout_rsci_ivld_run_sct(dout_rsci_ivld_run_sct)
    );
  decimator_run_dout_rsci_dout_wait_dp decimator_run_dout_rsci_dout_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run_din_rsci
// ------------------------------------------------------------------


module decimator_run_din_rsci (
  clk, rst, din_rsc_dat, din_rsc_vld, din_rsc_rdy, run_wen, din_rsci_oswt, din_rsci_wen_comp,
      din_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [7:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [7:0] din_rsci_idat_mxwt;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_bcwt;
  wire din_rsci_irdy_run_sct;
  wire din_rsci_ivld;
  wire [7:0] din_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd5),
  .width(32'sd8)) din_rsci (
      .rdy(din_rsc_rdy),
      .vld(din_rsc_vld),
      .dat(din_rsc_dat),
      .irdy(din_rsci_irdy_run_sct),
      .ivld(din_rsci_ivld),
      .idat(din_rsci_idat)
    );
  decimator_run_din_rsci_din_wait_ctrl decimator_run_din_rsci_din_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_irdy_run_sct(din_rsci_irdy_run_sct),
      .din_rsci_ivld(din_rsci_ivld)
    );
  decimator_run_din_rsci_din_wait_dp decimator_run_din_rsci_din_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_idat(din_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_run
// ------------------------------------------------------------------


module fir_run (
  clk, rst, input_rsc_dat, input_rsc_vld, input_rsc_rdy, coeffs, output_rsc_dat,
      output_rsc_vld, output_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [63:0] coeffs;
  output [7:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire input_rsci_wen_comp;
  wire [7:0] input_rsci_idat_mxwt;
  wire output_rsci_wen_comp;
  reg [7:0] output_rsci_idat;
  wire [9:0] fsm_output;
  wire or_22_tmp;
  wire MAC_and_4_ssc;
  reg reg_output_rsci_iswt0_cse;
  reg reg_input_rsci_iswt0_cse;
  wire MAC_and_cse;
  reg [7:0] reg_MAC_asn_8_cse;
  reg [7:0] reg_MAC_asn_4_cse;
  wire MAC_acc_8_itm_mx0c0;
  wire MAC_acc_8_itm_mx0c1;
  wire [15:0] z_out;
  wire [16:0] z_out_1;
  wire [17:0] nl_z_out_1;
  wire [17:0] z_out_2;
  wire [18:0] nl_z_out_2;
  reg [7:0] regs_2_sva;
  reg [7:0] regs_6_sva;
  reg [7:0] regs_0_sva;
  reg [15:0] MAC_3_mul_itm;
  reg [7:0] MAC_asn_10_itm;
  reg [7:0] MAC_asn_12_itm;
  reg [16:0] MAC_acc_7_itm;
  reg MAC_acc_8_itm_17;
  reg [8:0] MAC_acc_8_itm_16_8;
  reg [7:0] MAC_acc_8_itm_7_0;

  wire[18:0] MAC_8_acc_1_nl;
  wire[19:0] nl_MAC_8_acc_1_nl;
  wire MAC_and_8_nl;
  wire MAC_and_6_nl;
  wire[7:0] MAC_mux1h_6_nl;
  wire[7:0] MAC_mux1h_7_nl;
  wire signed [15:0] nl_mul_sgnd;
  wire[15:0] MAC_mux_6_nl;
  wire[15:0] MAC_MAC_mux_2_nl;
  wire[8:0] MAC_mux_7_nl;
  wire[7:0] MAC_mux_8_nl;
  wire[16:0] MAC_mux_9_nl;

  // Interconnect Declarations for Component Instantiations 
  fir_run_input_rsci fir_run_input_rsci_inst (
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .input_rsci_oswt(reg_input_rsci_iswt0_cse),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .input_rsci_idat_mxwt(input_rsci_idat_mxwt)
    );
  fir_run_output_rsci fir_run_output_rsci_inst (
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .output_rsci_oswt(reg_output_rsci_iswt0_cse),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_idat(output_rsci_idat)
    );
  fir_run_staller fir_run_staller_inst (
      .run_wen(run_wen),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .output_rsci_wen_comp(output_rsci_wen_comp)
    );
  fir_run_run_fsm fir_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign MAC_and_cse = run_wen & (fsm_output[9]);
  assign or_22_tmp = (fsm_output[3:2]!=2'b00);
  assign MAC_and_4_ssc = run_wen & (MAC_acc_8_itm_mx0c0 | MAC_acc_8_itm_mx0c1 | (fsm_output[6]));
  assign MAC_acc_8_itm_mx0c0 = (fsm_output[3:1]!=3'b000);
  assign MAC_acc_8_itm_mx0c1 = (fsm_output[5:4]!=2'b00);
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_idat <= 8'b00000000;
    end
    else if ( run_wen & (fsm_output[8]) ) begin
      output_rsci_idat <= readslicef_19_8_11(MAC_8_acc_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_output_rsci_iswt0_cse <= 1'b0;
      reg_input_rsci_iswt0_cse <= 1'b0;
      MAC_3_mul_itm <= 16'b0000000000000000;
    end
    else if ( run_wen ) begin
      reg_output_rsci_iswt0_cse <= fsm_output[8];
      reg_input_rsci_iswt0_cse <= (fsm_output[0]) | (fsm_output[9]);
      MAC_3_mul_itm <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_asn_10_itm <= 8'b00000000;
      reg_MAC_asn_8_cse <= 8'b00000000;
      regs_2_sva <= 8'b00000000;
      reg_MAC_asn_4_cse <= 8'b00000000;
      regs_6_sva <= 8'b00000000;
    end
    else if ( MAC_and_cse ) begin
      MAC_asn_10_itm <= reg_MAC_asn_4_cse;
      reg_MAC_asn_8_cse <= MAC_asn_10_itm;
      regs_2_sva <= MAC_asn_12_itm;
      reg_MAC_asn_4_cse <= regs_2_sva;
      regs_6_sva <= reg_MAC_asn_8_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_0_sva <= 8'b00000000;
    end
    else if ( run_wen & (fsm_output[4]) ) begin
      regs_0_sva <= MAC_acc_8_itm_7_0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_asn_12_itm <= 8'b00000000;
    end
    else if ( run_wen & ((fsm_output[9]) | (fsm_output[3])) ) begin
      MAC_asn_12_itm <= MUX_v_8_2_2(regs_0_sva, regs_6_sva, fsm_output[9]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_8_itm_17 <= 1'b0;
    end
    else if ( MAC_and_4_ssc ) begin
      MAC_acc_8_itm_17 <= z_out_2[17];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_8_itm_16_8 <= 9'b000000000;
    end
    else if ( MAC_and_4_ssc & (~ (fsm_output[5])) ) begin
      MAC_acc_8_itm_16_8 <= MUX_v_9_2_2((z_out_1[16:8]), (z_out_2[16:8]), fsm_output[6]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_8_itm_7_0 <= 8'b00000000;
    end
    else if ( MAC_and_4_ssc & (~(or_22_tmp | (fsm_output[5]))) ) begin
      MAC_acc_8_itm_7_0 <= MUX1HOT_v_8_3_2(input_rsci_idat_mxwt, (z_out_1[7:0]),
          (z_out_2[7:0]), {MAC_and_8_nl , MAC_and_6_nl , (fsm_output[6])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_7_itm <= 17'b00000000000000000;
    end
    else if ( run_wen & (fsm_output[2]) ) begin
      MAC_acc_7_itm <= z_out_1;
    end
  end
  assign nl_MAC_8_acc_1_nl = conv_s2s_18_19({MAC_acc_8_itm_17 , MAC_acc_8_itm_16_8
      , MAC_acc_8_itm_7_0}) + conv_s2s_18_19(z_out_2);
  assign MAC_8_acc_1_nl = nl_MAC_8_acc_1_nl[18:0];
  assign MAC_and_8_nl = (~ or_22_tmp) & MAC_acc_8_itm_mx0c0;
  assign MAC_and_6_nl = (~ (fsm_output[5])) & MAC_acc_8_itm_mx0c1;
  assign MAC_mux1h_6_nl = MUX1HOT_v_8_8_2((coeffs[39:32]), (coeffs[55:48]), (coeffs[15:8]),
      (coeffs[31:24]), (coeffs[47:40]), (coeffs[7:0]), (coeffs[23:16]), (coeffs[63:56]),
      {(fsm_output[8]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[2])});
  assign MAC_mux1h_7_nl = MUX1HOT_v_8_8_2(MAC_asn_10_itm, regs_6_sva, regs_0_sva,
      reg_MAC_asn_4_cse, reg_MAC_asn_8_cse, MAC_acc_8_itm_7_0, regs_2_sva, MAC_asn_12_itm,
      {(fsm_output[8]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[2])});
  assign nl_mul_sgnd = $signed(MAC_mux1h_6_nl) * $signed(MAC_mux1h_7_nl);
  assign z_out = $unsigned(nl_mul_sgnd);
  assign MAC_mux_6_nl = MUX_v_16_2_2(MAC_3_mul_itm, z_out, fsm_output[2]);
  assign MAC_MAC_mux_2_nl = MUX_v_16_2_2(z_out, MAC_3_mul_itm, fsm_output[2]);
  assign nl_z_out_1 = conv_s2u_16_17(MAC_mux_6_nl) + conv_s2u_16_17(MAC_MAC_mux_2_nl);
  assign z_out_1 = nl_z_out_1[16:0];
  assign MAC_mux_7_nl = MUX_v_9_2_2((z_out_1[16:8]), MAC_acc_8_itm_16_8, fsm_output[6]);
  assign MAC_mux_8_nl = MUX_v_8_2_2((z_out_1[7:0]), MAC_acc_8_itm_7_0, fsm_output[6]);
  assign MAC_mux_9_nl = MUX_v_17_2_2(MAC_acc_7_itm, z_out_1, fsm_output[6]);
  assign nl_z_out_2 = conv_s2u_17_18({MAC_mux_7_nl , MAC_mux_8_nl}) + conv_s2u_17_18(MAC_mux_9_nl);
  assign z_out_2 = nl_z_out_2[17:0];

  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_8_2;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [7:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    MUX1HOT_v_8_8_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input  sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [7:0] readslicef_19_8_11;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_19_8_11 = tmp[7:0];
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [16:0] conv_s2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator_run
// ------------------------------------------------------------------


module decimator_run (
  clk, rst, din_rsc_dat, din_rsc_vld, din_rsc_rdy, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  output [7:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire din_rsci_wen_comp;
  wire [7:0] din_rsci_idat_mxwt;
  wire dout_rsci_wen_comp;
  reg [7:0] dout_rsci_idat;
  wire [1:0] fsm_output;
  wire equal_tmp;
  reg reg_dout_rsci_iswt0_cse;
  reg reg_din_rsci_iswt0_cse;
  reg [1:0] count_2_0_sva_1_0;
  wire [2:0] nl_count_2_0_sva_1_0;


  // Interconnect Declarations for Component Instantiations 
  decimator_run_din_rsci decimator_run_din_rsci_inst (
      .clk(clk),
      .rst(rst),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .run_wen(run_wen),
      .din_rsci_oswt(reg_din_rsci_iswt0_cse),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt)
    );
  decimator_run_dout_rsci decimator_run_dout_rsci_inst (
      .clk(clk),
      .rst(rst),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .run_wen(run_wen),
      .dout_rsci_oswt(reg_dout_rsci_iswt0_cse),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_idat(dout_rsci_idat)
    );
  decimator_run_staller decimator_run_staller_inst (
      .run_wen(run_wen),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .dout_rsci_wen_comp(dout_rsci_wen_comp)
    );
  decimator_run_run_fsm decimator_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign equal_tmp = ~((count_2_0_sva_1_0!=2'b00));
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_idat <= 8'b00000000;
    end
    else if ( run_wen & (~((~ equal_tmp) | (fsm_output[0]))) ) begin
      dout_rsci_idat <= din_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_dout_rsci_iswt0_cse <= 1'b0;
      reg_din_rsci_iswt0_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_dout_rsci_iswt0_cse <= equal_tmp & (fsm_output[1]);
      reg_din_rsci_iswt0_cse <= 1'b1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      count_2_0_sva_1_0 <= 2'b00;
    end
    else if ( run_wen & (~ (fsm_output[0])) ) begin
      count_2_0_sva_1_0 <= nl_count_2_0_sva_1_0[1:0];
    end
  end
  assign nl_count_2_0_sva_1_0  = count_2_0_sva_1_0 + 2'b01;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, input_rsc_dat, input_rsc_vld, input_rsc_rdy, coeffs, output_rsc_dat,
      output_rsc_vld, output_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [63:0] coeffs;
  output [7:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  fir_run fir_run_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .coeffs(coeffs),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    decimator
// ------------------------------------------------------------------


module decimator (
  clk, rst, din_rsc_dat, din_rsc_vld, din_rsc_rdy, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  output [7:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  decimator_run decimator_run_inst (
      .clk(clk),
      .rst(rst),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    top
// ------------------------------------------------------------------


module top (
  clk, rst, din_rsc_dat, din_rsc_vld, din_rsc_rdy, coeffs, dout_rsc_dat, dout_rsc_vld,
      dout_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input [63:0] coeffs;
  output [7:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;


  // Interconnect Declarations
  wire [7:0] output_rsc_dat_n_block0;
  wire [7:0] output_rsc_dat_n_block1;
  wire [7:0] dout_rsc_dat_n_block2;
  wire input_rsc_rdy_n_block0_bud;
  wire output_rsc_vld_n_block0_bud;
  wire input_rsc_rdy_n_block1_bud;
  wire output_rsc_vld_n_block1_bud;
  wire din_rsc_rdy_n_block2_bud;
  wire dout_rsc_vld_n_block2_bud;


  // Interconnect Declarations for Component Instantiations 
  fir block0 (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(din_rsc_dat),
      .input_rsc_vld(din_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy_n_block0_bud),
      .coeffs(coeffs),
      .output_rsc_dat(output_rsc_dat_n_block0),
      .output_rsc_vld(output_rsc_vld_n_block0_bud),
      .output_rsc_rdy(input_rsc_rdy_n_block1_bud)
    );
  fir block1 (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(output_rsc_dat_n_block0),
      .input_rsc_vld(output_rsc_vld_n_block0_bud),
      .input_rsc_rdy(input_rsc_rdy_n_block1_bud),
      .coeffs(coeffs),
      .output_rsc_dat(output_rsc_dat_n_block1),
      .output_rsc_vld(output_rsc_vld_n_block1_bud),
      .output_rsc_rdy(din_rsc_rdy_n_block2_bud)
    );
  decimator block2 (
      .clk(clk),
      .rst(rst),
      .din_rsc_dat(output_rsc_dat_n_block1),
      .din_rsc_vld(output_rsc_vld_n_block1_bud),
      .din_rsc_rdy(din_rsc_rdy_n_block2_bud),
      .dout_rsc_dat(dout_rsc_dat_n_block2),
      .dout_rsc_vld(dout_rsc_vld_n_block2_bud),
      .dout_rsc_rdy(dout_rsc_rdy)
    );
  assign din_rsc_rdy = input_rsc_rdy_n_block0_bud;
  assign dout_rsc_vld = dout_rsc_vld_n_block2_bud;
  assign dout_rsc_dat = dout_rsc_dat_n_block2;
endmodule



